/*
	Okay, actually I'm going to build something more interesting.
	I want to build a verilog SAT solver
*/



module myModule();

initial
  begin
    $display("Hello World!");
    $finish ;
  end

endmodule
